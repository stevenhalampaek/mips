/************************************************************
 * Author: 
 * Description:
 ************************************************************/

module ();

endmodule
